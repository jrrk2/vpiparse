module logand (
    input [1:0] a,
    input [1:0] b,
    output y);

    assign
      y = a && b;

endmodule
