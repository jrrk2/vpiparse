module op_priority(input [3:0] u1, u2, u3, output [3:0] y);

   assign y = u1 + u2 * u3;

endmodule
