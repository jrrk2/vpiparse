module mult(
    output wire [3:0] out1,
    input wire [3:0] arg1);
   
   assign out1 = arg1;

endmodule

module add(
    output wire [3:0] out1,
    input wire [3:0] arg1);
   
   assign out1 = arg1;

endmodule
	   
