module index;

   wire [7:0] data;

   assign data[7:0] = 8'b1;

endmodule // index
