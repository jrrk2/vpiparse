module equal(input [3:0] u1, u2, output y);

   assign y = u1 == u2;

endmodule
