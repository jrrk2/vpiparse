module one;
	wire x;
endmodule
module three;
	wire x;
endmodule
module two;
	wire x;
endmodule